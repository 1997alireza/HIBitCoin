library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package sha_functions is
end sha_functions;

package body sha_functions is

end package body;